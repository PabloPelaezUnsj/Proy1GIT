library ieee;
use ieee.std_logic_1164.all;

entity Proy1GIT is
			port(	x1, x2: in	std_logic_vector(3 downto 0);
					displays: out std_logic_vector(13 downto 0) );
end Proy1GIT;


architecture bev of Proy1GIT

begin

--TODO




end bev;

	